// vidor_sys.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module vidor_sys (
		input  wire       clk_clk,                                                    //                      clk.clk
		input  wire       myocontrol_0_conduit_end_angle_miso,                        // myocontrol_0_conduit_end.angle_miso
		output wire       myocontrol_0_conduit_end_angle_mosi,                        //                         .angle_mosi
		output wire       myocontrol_0_conduit_end_angle_sck,                         //                         .angle_sck
		output wire [3:0] myocontrol_0_conduit_end_angle_ss_n_o,                      //                         .angle_ss_n_o
		output wire       myocontrol_0_conduit_end_gpio_n,                            //                         .gpio_n
		input  wire       myocontrol_0_conduit_end_mirrored_muscle_unit,              //                         .mirrored_muscle_unit
		input  wire       myocontrol_0_conduit_end_miso,                              //                         .miso
		output wire       myocontrol_0_conduit_end_mosi,                              //                         .mosi
		input  wire       myocontrol_0_conduit_end_power_sense_n,                     //                         .power_sense_n
		output wire [3:0] myocontrol_0_conduit_end_ss_n_o,                            //                         .ss_n_o
		output wire       myocontrol_0_conduit_end_sck,                               //                         .sck
		input  wire       reset_reset_n,                                              //                    reset.reset_n
		input  wire       spi_bridge_mosi_to_the_spislave_inst_for_spichain,          //               spi_bridge.mosi_to_the_spislave_inst_for_spichain
		input  wire       spi_bridge_nss_to_the_spislave_inst_for_spichain,           //                         .nss_to_the_spislave_inst_for_spichain
		inout  wire       spi_bridge_miso_to_and_from_the_spislave_inst_for_spichain, //                         .miso_to_and_from_the_spislave_inst_for_spichain
		input  wire       spi_bridge_sclk_to_the_spislave_inst_for_spichain           //                         .sclk_to_the_spislave_inst_for_spichain
	);

	wire  [31:0] spi_avalon_bridge_avalon_master_readdata;                  // mm_interconnect_0:spi_avalon_bridge_avalon_master_readdata -> spi_avalon_bridge:readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire         spi_avalon_bridge_avalon_master_waitrequest;               // mm_interconnect_0:spi_avalon_bridge_avalon_master_waitrequest -> spi_avalon_bridge:waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire  [31:0] spi_avalon_bridge_avalon_master_address;                   // spi_avalon_bridge:address_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_avalon_bridge_avalon_master_address
	wire   [3:0] spi_avalon_bridge_avalon_master_byteenable;                // spi_avalon_bridge:byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_avalon_bridge_avalon_master_byteenable
	wire         spi_avalon_bridge_avalon_master_read;                      // spi_avalon_bridge:read_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_avalon_bridge_avalon_master_read
	wire         spi_avalon_bridge_avalon_master_readdatavalid;             // mm_interconnect_0:spi_avalon_bridge_avalon_master_readdatavalid -> spi_avalon_bridge:readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain
	wire         spi_avalon_bridge_avalon_master_write;                     // spi_avalon_bridge:write_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_avalon_bridge_avalon_master_write
	wire  [31:0] spi_avalon_bridge_avalon_master_writedata;                 // spi_avalon_bridge:writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:spi_avalon_bridge_avalon_master_writedata
	wire  [31:0] mm_interconnect_0_myocontrol_0_avalon_slave_0_readdata;    // MYOControl_0:readdata -> mm_interconnect_0:MYOControl_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_myocontrol_0_avalon_slave_0_waitrequest; // MYOControl_0:waitrequest -> mm_interconnect_0:MYOControl_0_avalon_slave_0_waitrequest
	wire  [15:0] mm_interconnect_0_myocontrol_0_avalon_slave_0_address;     // mm_interconnect_0:MYOControl_0_avalon_slave_0_address -> MYOControl_0:address
	wire         mm_interconnect_0_myocontrol_0_avalon_slave_0_read;        // mm_interconnect_0:MYOControl_0_avalon_slave_0_read -> MYOControl_0:read
	wire         mm_interconnect_0_myocontrol_0_avalon_slave_0_write;       // mm_interconnect_0:MYOControl_0_avalon_slave_0_write -> MYOControl_0:write
	wire  [31:0] mm_interconnect_0_myocontrol_0_avalon_slave_0_writedata;   // mm_interconnect_0:MYOControl_0_avalon_slave_0_writedata -> MYOControl_0:writedata
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [MYOControl_0:reset, mm_interconnect_0:spi_avalon_bridge_clk_reset_reset_bridge_in_reset_reset, spi_avalon_bridge:reset_n]

	MYOControl #(
		.NUMBER_OF_MOTORS        (4),
		.CLOCK_SPEED_HZ          (24000000),
		.ENABLE_MYOBRICK_CONTROL (0)
	) myocontrol_0 (
		.reset                (rst_controller_reset_out_reset),                            //          reset.reset
		.address              (mm_interconnect_0_myocontrol_0_avalon_slave_0_address),     // avalon_slave_0.address
		.write                (mm_interconnect_0_myocontrol_0_avalon_slave_0_write),       //               .write
		.writedata            (mm_interconnect_0_myocontrol_0_avalon_slave_0_writedata),   //               .writedata
		.read                 (mm_interconnect_0_myocontrol_0_avalon_slave_0_read),        //               .read
		.readdata             (mm_interconnect_0_myocontrol_0_avalon_slave_0_readdata),    //               .readdata
		.waitrequest          (mm_interconnect_0_myocontrol_0_avalon_slave_0_waitrequest), //               .waitrequest
		.angle_miso           (myocontrol_0_conduit_end_angle_miso),                       //    conduit_end.angle_miso
		.angle_mosi           (myocontrol_0_conduit_end_angle_mosi),                       //               .angle_mosi
		.angle_sck            (myocontrol_0_conduit_end_angle_sck),                        //               .angle_sck
		.angle_ss_n_o         (myocontrol_0_conduit_end_angle_ss_n_o),                     //               .angle_ss_n_o
		.gpio_n               (myocontrol_0_conduit_end_gpio_n),                           //               .gpio_n
		.mirrored_muscle_unit (myocontrol_0_conduit_end_mirrored_muscle_unit),             //               .mirrored_muscle_unit
		.miso                 (myocontrol_0_conduit_end_miso),                             //               .miso
		.mosi                 (myocontrol_0_conduit_end_mosi),                             //               .mosi
		.power_sense_n        (myocontrol_0_conduit_end_power_sense_n),                    //               .power_sense_n
		.ss_n_o               (myocontrol_0_conduit_end_ss_n_o),                           //               .ss_n_o
		.sck                  (myocontrol_0_conduit_end_sck),                              //               .sck
		.clock                (clk_clk)                                                    //     clock_sink.clk
	);

	SPISlaveToAvalonMasterBridge #(
		.SYNC_DEPTH (5)
	) spi_avalon_bridge (
		.clk                                                                    (clk_clk),                                                    //           clk.clk
		.reset_n                                                                (~rst_controller_reset_out_reset),                            //     clk_reset.reset_n
		.mosi_to_the_spislave_inst_for_spichain                                 (spi_bridge_mosi_to_the_spislave_inst_for_spichain),          //      export_0.export
		.nss_to_the_spislave_inst_for_spichain                                  (spi_bridge_nss_to_the_spislave_inst_for_spichain),           //              .export
		.miso_to_and_from_the_spislave_inst_for_spichain                        (spi_bridge_miso_to_and_from_the_spislave_inst_for_spichain), //              .export
		.sclk_to_the_spislave_inst_for_spichain                                 (spi_bridge_sclk_to_the_spislave_inst_for_spichain),          //              .export
		.address_from_the_altera_avalon_packets_to_master_inst_for_spichain     (spi_avalon_bridge_avalon_master_address),                    // avalon_master.address
		.byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain  (spi_avalon_bridge_avalon_master_byteenable),                 //              .byteenable
		.read_from_the_altera_avalon_packets_to_master_inst_for_spichain        (spi_avalon_bridge_avalon_master_read),                       //              .read
		.readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain      (spi_avalon_bridge_avalon_master_readdata),                   //              .readdata
		.readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain (spi_avalon_bridge_avalon_master_readdatavalid),              //              .readdatavalid
		.waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain   (spi_avalon_bridge_avalon_master_waitrequest),                //              .waitrequest
		.write_from_the_altera_avalon_packets_to_master_inst_for_spichain       (spi_avalon_bridge_avalon_master_write),                      //              .write
		.writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain   (spi_avalon_bridge_avalon_master_writedata)                   //              .writedata
	);

	vidor_sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                           (clk_clk),                                                   //                                         clk_0_clk.clk
		.spi_avalon_bridge_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // spi_avalon_bridge_clk_reset_reset_bridge_in_reset.reset
		.spi_avalon_bridge_avalon_master_address                 (spi_avalon_bridge_avalon_master_address),                   //                   spi_avalon_bridge_avalon_master.address
		.spi_avalon_bridge_avalon_master_waitrequest             (spi_avalon_bridge_avalon_master_waitrequest),               //                                                  .waitrequest
		.spi_avalon_bridge_avalon_master_byteenable              (spi_avalon_bridge_avalon_master_byteenable),                //                                                  .byteenable
		.spi_avalon_bridge_avalon_master_read                    (spi_avalon_bridge_avalon_master_read),                      //                                                  .read
		.spi_avalon_bridge_avalon_master_readdata                (spi_avalon_bridge_avalon_master_readdata),                  //                                                  .readdata
		.spi_avalon_bridge_avalon_master_readdatavalid           (spi_avalon_bridge_avalon_master_readdatavalid),             //                                                  .readdatavalid
		.spi_avalon_bridge_avalon_master_write                   (spi_avalon_bridge_avalon_master_write),                     //                                                  .write
		.spi_avalon_bridge_avalon_master_writedata               (spi_avalon_bridge_avalon_master_writedata),                 //                                                  .writedata
		.MYOControl_0_avalon_slave_0_address                     (mm_interconnect_0_myocontrol_0_avalon_slave_0_address),     //                       MYOControl_0_avalon_slave_0.address
		.MYOControl_0_avalon_slave_0_write                       (mm_interconnect_0_myocontrol_0_avalon_slave_0_write),       //                                                  .write
		.MYOControl_0_avalon_slave_0_read                        (mm_interconnect_0_myocontrol_0_avalon_slave_0_read),        //                                                  .read
		.MYOControl_0_avalon_slave_0_readdata                    (mm_interconnect_0_myocontrol_0_avalon_slave_0_readdata),    //                                                  .readdata
		.MYOControl_0_avalon_slave_0_writedata                   (mm_interconnect_0_myocontrol_0_avalon_slave_0_writedata),   //                                                  .writedata
		.MYOControl_0_avalon_slave_0_waitrequest                 (mm_interconnect_0_myocontrol_0_avalon_slave_0_waitrequest)  //                                                  .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
